Spice circuit Gen

R1 w2 0 5
R2D2 w1 0 4
V w2 w1 10
.options savecurrents

.control
op
print V(w1)
print V(w2)
print @R1[i]
print @R2D2[i]
print I(V)
exit
.endc
.end
