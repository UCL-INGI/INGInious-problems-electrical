Spice circuit Gen

R1 0 w1 5
R2D2 0 w0 4
V w0 w1 10
.options savecurrents

.control
op
print V(w0)
print V(w1)
print @R1[i]
print @R2D2[i]
print I(V)
exit
.endc
.end
