Spice circuit Gen

R1 0 w1 5
V2 0 w2 5
V w1 w2 10
.options savecurrents

.control
op
print V(w1)
print V(w2)
print @R1[i]
print I(V2)
print I(V)
exit
.endc
.end
