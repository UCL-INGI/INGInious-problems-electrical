Spice circuit Gen

R1 w0 0 5
V w0 0 10
.options savecurrents

.control
op
print V(w0)
print @R1[i]
print I(V)
exit
.endc
.end
